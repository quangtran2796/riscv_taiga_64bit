package Taiga;

interface Taiga;
// Add custom interface definitions
endinterface

module mkTaiga(Taiga);

    rule doNothing;
        $display("Hello World!");
    endrule

endmodule

endpackage
